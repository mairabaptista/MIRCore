module BIOS(address, biosOut, clk_auto);

	input [31:0]address;
	input clk_auto;
	output reg [31:0]biosOut;
	
	reg [31:0] bios[63:0];
	initial
		begin				
bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000100; // addi: $sp = $sp + (4)
bios[2] <= 32'b001111_00000_10100_0000000000000001; // li: load 1 in register $t0
bios[3] <= 32'b010000_11110_10100_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t0]
bios[4] <= 32'b001111_00000_10101_0110000110101000; // li: load 25000 in register $t1
bios[5] <= 32'b010000_11110_10101_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t1]
bios[6] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[7] <= 32'b001111_00000_10110_0000000000001010; // li: load 10 in register $t2
bios[8] <= 32'b110000_01010_10110_10111_00000000000; // lt: if($s0 < $t2): $t3 = 1, else $t3 = 0
bios[9] <= 32'b010001_10111_00000_0000000000010010; // bneq: if($t3 == 0) jump to 18
bios[10] <= 32'b001110_11110_01011_1111111111111110; // lw: $s1 = mem[$sp] + (-2)
bios[11] <= 32'b001100_01011_11000_0110000110101000; // addi: $t4 = $s1 + (25000)
bios[12] <= 32'b010000_11110_11000_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t4]
bios[13] <= 32'b001110_11110_01011_1111111111111110; // lw: $s1 = mem[$sp] + (-2)
bios[14] <= 32'b001100_01010_11001_0000000000000001; // addi: $t5 = $s0 + (1)
bios[15] <= 32'b010000_11110_11001_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t5]
bios[16] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[17] <= 32'b011010_00000000000000000000000110; // jump to 6 (L1)
bios[18] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
bios[19] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[20] <= 32'b101101_00000_00110_0000000000000000; // baud $a0
bios[21] <= 32'b011100_00000000000000000000000000; // nop
bios[22] <= 32'b101111_00000_11010_0000000000000000; // rcv $t6
bios[23] <= 32'b010000_11110_11010_0000000000000000; // sw: mem[$sp + (0)] = mem[$t6]
bios[24] <= 32'b001110_11110_01011_0000000000000000; // lw: $s1 = mem[$sp] + (0)
bios[25] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
bios[26] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[27] <= 32'b001101_11110_11110_0000000000000100; // subi: $sp = $sp - (4)
bios[28] <= 32'b011101_00000000000000000000000000; // hlt

/*bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000101; // addi: $sp = $sp + (5)
bios[2] <= 32'b001111_00000_00110_0000000000001010; // li: load 10 in register $a0
bios[3] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
bios[4] <= 32'b011100_00000000000000000000000000; // nop
bios[5] <= 32'b100101_00000_10100_0000000000000000; // in $t0
bios[6] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
bios[7] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
bios[8] <= 32'b001100_01010_10101_0000000000000010; // addi: $t1 = $s0 + (2)
bios[9] <= 32'b010000_11110_10101_0000000000000000; // sw: mem[$sp + (0)] = mem[$t1]
bios[10] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
bios[11] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[12] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[13] <= 32'b001111_00000_10110_0000000000000000; // li: load 0 in register $t2
bios[14] <= 32'b010000_11110_10110_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t2]
bios[15] <= 32'b001110_11110_01010_1111111111111101; // lw: $s0 = mem[$sp] + (-3)
bios[16] <= 32'b001111_00000_10111_0000010000000000; // li: load 1024 in register $t3
bios[17] <= 32'b100010_01010_10111_11000_00000000000; // neq: if($s0 != $t3): $t4 = 1, else $t4 = 0
bios[18] <= 32'b010001_11000_00000_0000000000011110; // bneq: if($t4 == 0) jump to 30
bios[19] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[20] <= 32'b110010_00110_11001_0000000000000000; // lhd: $t5 = hd[$a0]
bios[21] <= 32'b010000_11110_11001_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t5]
bios[22] <= 32'b001110_11110_01011_1111111111111110; // lw: $s1 = mem[$sp] + (-2)
bios[23] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
bios[24] <= 32'b011011_01010_00111_0000000000000000; // mov: $a1 = $s0
bios[25] <= 32'b110101_00111_00110_0000000000000000; // smem: mem[$a0] = $a1
bios[26] <= 32'b001100_01010_11010_0000000000000001; // addi: $t6 = $s0 + (1)
bios[27] <= 32'b010000_11110_11010_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t6]
bios[28] <= 32'b001110_11110_01010_1111111111111101; // lw: $s0 = mem[$sp] + (-3)
bios[29] <= 32'b011010_00000000000000000000001111; // jump to 15 (L1)
bios[30] <= 32'b001111_00000_00110_0000000000001011; // li: load 11 in register $a0
bios[31] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
bios[32] <= 32'b011100_00000000000000000000000000; // nop
bios[33] <= 32'b100101_00000_11011_0000000000000000; // in $t7
bios[34] <= 32'b010000_11110_11011_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t7]
bios[35] <= 32'b001101_11110_11110_0000000000000101; // subi: $sp = $sp - (5)
bios[36] <= 32'b011101_00000000000000000000000000; // hlt*/





		end
	
	always @(posedge clk_auto)
		begin
			biosOut <= bios[address];
		end

	
endmodule

