module HD(clk_auto, clk, write_flag, input_data, hd_output, address) ;

	parameter DATA_WIDTH = 32; 
	parameter ADDR_WIDTH = 15; 
	parameter MAX_PROC_NUM = 16; 
	parameter REGION = (2**ADDR_WIDTH)/MAX_PROC_NUM;// 2048
	parameter DISK_SIZE = 4096;
	
	//INPUTS
	input clk_auto, clk, write_flag; //precisa do clk_auto?
	input [(DATA_WIDTH-1):0] input_data;  //data in -> to disk
	input [(DATA_WIDTH-1):0] address; //disk address
	
	//OUTPUTS
	output reg [(DATA_WIDTH-1):0] hd_output; //data out -> from disk 
	
	reg[(DATA_WIDTH-1):0] hd[DISK_SIZE-1:0]; //disk cells
	
	initial
	begin
	//OS
hd[0] <= 32'b011010_00000000000000001100101010; // jump to 810 (main)
hd[1] <= 32'b001100_11110_11110_0000000000000100; // addi: $sp = $sp + (4)
hd[2] <= 32'b010000_11110_00110_1111111111111111; // sw: mem[$sp + (-1)] = mem[$a0]
hd[3] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[4] <= 32'b001100_01010_10100_0000000000000001; // addi: $t0 = $s0 + (1)
hd[5] <= 32'b010000_11110_10100_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t0]
hd[6] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[7] <= 32'b001110_00101_01011_0000000000000001; // lw: $s1 = mem[$gp] + (1)
hd[8] <= 32'b000111_01010_01011_10101_00000000000; // mul: $t1 = $s0 * $s1
hd[9] <= 32'b010000_11110_10101_0000000000000000; // sw: mem[$sp + (0)] = mem[$t1]
hd[10] <= 32'b001111_00000_00110_0000000000000001; // li: load 1 in register $a0
hd[11] <= 32'b001110_11110_01100_0000000000000000; // lw: $s2 = mem[$sp] + (0)
hd[12] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[13] <= 32'b001111_00000_01000_0000000000000001; // li: load 1 in register $a2
hd[14] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[15] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[16] <= 32'b011011_00001_00110_0000000000000000; // mov: $a0 = $v0
hd[17] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[18] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[19] <= 32'b001111_00000_00110_0000000000000010; // li: load 2 in register $a0
hd[20] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[21] <= 32'b001111_00000_01000_0000000000000010; // li: load 2 in register $a2
hd[22] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[23] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[24] <= 32'b011011_00010_00110_0000000000000000; // mov: $a0 = $v1
hd[25] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[26] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[27] <= 32'b001111_00000_00110_0000000000000011; // li: load 3 in register $a0
hd[28] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[29] <= 32'b001111_00000_01000_0000000000000011; // li: load 3 in register $a2
hd[30] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[31] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[32] <= 32'b011011_00011_00110_0000000000000000; // mov: $a0 = $out1
hd[33] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[34] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[35] <= 32'b001111_00000_00110_0000000000000100; // li: load 4 in register $a0
hd[36] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[37] <= 32'b001111_00000_01000_0000000000000100; // li: load 4 in register $a2
hd[38] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[39] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[40] <= 32'b011011_00100_00110_0000000000000000; // mov: $a0 = $out2
hd[41] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[42] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[43] <= 32'b001111_00000_00110_0000000000000101; // li: load 5 in register $a0
hd[44] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[45] <= 32'b001111_00000_01000_0000000000000101; // li: load 5 in register $a2
hd[46] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[47] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[48] <= 32'b011011_00101_00110_0000000000000000; // mov: $a0 = $gp
hd[49] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[50] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[51] <= 32'b001111_00000_00110_0000000000000110; // li: load 6 in register $a0
hd[52] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[53] <= 32'b001111_00000_01000_0000000000000110; // li: load 6 in register $a2
hd[54] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[55] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[56] <= 32'b011011_00110_00110_0000000000000000; // mov: $a0 = $a0
hd[57] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[58] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[59] <= 32'b001111_00000_00110_0000000000000111; // li: load 7 in register $a0
hd[60] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[61] <= 32'b001111_00000_01000_0000000000000111; // li: load 7 in register $a2
hd[62] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[63] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[64] <= 32'b011011_00111_00110_0000000000000000; // mov: $a0 = $a1
hd[65] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[66] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[67] <= 32'b001111_00000_00110_0000000000001000; // li: load 8 in register $a0
hd[68] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[69] <= 32'b001111_00000_01000_0000000000001000; // li: load 8 in register $a2
hd[70] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[71] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[72] <= 32'b011011_01000_00110_0000000000000000; // mov: $a0 = $a2
hd[73] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[74] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[75] <= 32'b001111_00000_00110_0000000000001001; // li: load 9 in register $a0
hd[76] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[77] <= 32'b001111_00000_01000_0000000000001001; // li: load 9 in register $a2
hd[78] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[79] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[80] <= 32'b011011_01001_00110_0000000000000000; // mov: $a0 = $a3
hd[81] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[82] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[83] <= 32'b001111_00000_00110_0000000000001010; // li: load 10 in register $a0
hd[84] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[85] <= 32'b001111_00000_01000_0000000000001010; // li: load 10 in register $a2
hd[86] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[87] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[88] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[89] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[90] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[91] <= 32'b001111_00000_00110_0000000000001011; // li: load 11 in register $a0
hd[92] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[93] <= 32'b001111_00000_01000_0000000000001011; // li: load 11 in register $a2
hd[94] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[95] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[96] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
hd[97] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[98] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[99] <= 32'b001111_00000_00110_0000000000001100; // li: load 12 in register $a0
hd[100] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[101] <= 32'b001111_00000_01000_0000000000001100; // li: load 12 in register $a2
hd[102] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[103] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[104] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
hd[105] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[106] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[107] <= 32'b001111_00000_00110_0000000000001101; // li: load 13 in register $a0
hd[108] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[109] <= 32'b001111_00000_01000_0000000000001101; // li: load 13 in register $a2
hd[110] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[111] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[112] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
hd[113] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[114] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[115] <= 32'b001111_00000_00110_0000000000001110; // li: load 14 in register $a0
hd[116] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[117] <= 32'b001111_00000_01000_0000000000001110; // li: load 14 in register $a2
hd[118] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[119] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[120] <= 32'b011011_01110_00110_0000000000000000; // mov: $a0 = $s4
hd[121] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[122] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[123] <= 32'b001111_00000_00110_0000000000001111; // li: load 15 in register $a0
hd[124] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[125] <= 32'b001111_00000_01000_0000000000001111; // li: load 15 in register $a2
hd[126] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[127] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[128] <= 32'b011011_01111_00110_0000000000000000; // mov: $a0 = $s5
hd[129] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[130] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[131] <= 32'b001111_00000_00110_0000000000010000; // li: load 16 in register $a0
hd[132] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[133] <= 32'b001111_00000_01000_0000000000010000; // li: load 16 in register $a2
hd[134] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[135] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[136] <= 32'b011011_10000_00110_0000000000000000; // mov: $a0 = $s6
hd[137] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[138] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[139] <= 32'b001111_00000_00110_0000000000010001; // li: load 17 in register $a0
hd[140] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[141] <= 32'b001111_00000_01000_0000000000010001; // li: load 17 in register $a2
hd[142] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[143] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[144] <= 32'b011011_10001_00110_0000000000000000; // mov: $a0 = $s7
hd[145] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[146] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[147] <= 32'b001111_00000_00110_0000000000010010; // li: load 18 in register $a0
hd[148] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[149] <= 32'b001111_00000_01000_0000000000010010; // li: load 18 in register $a2
hd[150] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[151] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[152] <= 32'b011011_10010_00110_0000000000000000; // mov: $a0 = $s8
hd[153] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[154] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[155] <= 32'b001111_00000_00110_0000000000010011; // li: load 19 in register $a0
hd[156] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[157] <= 32'b001111_00000_01000_0000000000010011; // li: load 19 in register $a2
hd[158] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[159] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[160] <= 32'b011011_10011_00110_0000000000000000; // mov: $a0 = $s9
hd[161] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[162] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[163] <= 32'b001111_00000_00110_0000000000010100; // li: load 20 in register $a0
hd[164] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[165] <= 32'b001111_00000_01000_0000000000010100; // li: load 20 in register $a2
hd[166] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[167] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[168] <= 32'b011011_10100_00110_0000000000000000; // mov: $a0 = $t0
hd[169] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[170] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[171] <= 32'b001111_00000_00110_0000000000010101; // li: load 21 in register $a0
hd[172] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[173] <= 32'b001111_00000_01000_0000000000010101; // li: load 21 in register $a2
hd[174] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[175] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[176] <= 32'b011011_10101_00110_0000000000000000; // mov: $a0 = $t1
hd[177] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[178] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[179] <= 32'b001111_00000_00110_0000000000010110; // li: load 22 in register $a0
hd[180] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[181] <= 32'b001111_00000_01000_0000000000010110; // li: load 22 in register $a2
hd[182] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[183] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[184] <= 32'b011011_10110_00110_0000000000000000; // mov: $a0 = $t2
hd[185] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[186] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[187] <= 32'b001111_00000_00110_0000000000010111; // li: load 23 in register $a0
hd[188] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[189] <= 32'b001111_00000_01000_0000000000010111; // li: load 23 in register $a2
hd[190] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[191] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[192] <= 32'b011011_10111_00110_0000000000000000; // mov: $a0 = $t3
hd[193] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[194] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[195] <= 32'b001111_00000_00110_0000000000011000; // li: load 24 in register $a0
hd[196] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[197] <= 32'b001111_00000_01000_0000000000011000; // li: load 24 in register $a2
hd[198] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[199] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[200] <= 32'b011011_11000_00110_0000000000000000; // mov: $a0 = $t4
hd[201] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[202] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[203] <= 32'b001111_00000_00110_0000000000011001; // li: load 25 in register $a0
hd[204] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[205] <= 32'b001111_00000_01000_0000000000011001; // li: load 25 in register $a2
hd[206] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[207] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[208] <= 32'b011011_11001_00110_0000000000000000; // mov: $a0 = $t5
hd[209] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[210] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[211] <= 32'b001111_00000_00110_0000000000011010; // li: load 26 in register $a0
hd[212] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[213] <= 32'b001111_00000_01000_0000000000011010; // li: load 26 in register $a2
hd[214] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[215] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[216] <= 32'b011011_11010_00110_0000000000000000; // mov: $a0 = $t6
hd[217] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[218] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[219] <= 32'b001111_00000_00110_0000000000011011; // li: load 27 in register $a0
hd[220] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[221] <= 32'b001111_00000_01000_0000000000011011; // li: load 27 in register $a2
hd[222] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[223] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[224] <= 32'b011011_11011_00110_0000000000000000; // mov: $a0 = $t7
hd[225] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[226] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[227] <= 32'b001111_00000_00110_0000000000011100; // li: load 28 in register $a0
hd[228] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[229] <= 32'b001111_00000_01000_0000000000011100; // li: load 28 in register $a2
hd[230] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[231] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[232] <= 32'b011011_11100_00110_0000000000000000; // mov: $a0 = $t8
hd[233] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[234] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[235] <= 32'b001111_00000_00110_0000000000011101; // li: load 29 in register $a0
hd[236] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[237] <= 32'b001111_00000_01000_0000000000011101; // li: load 29 in register $a2
hd[238] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[239] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[240] <= 32'b011011_11101_00110_0000000000000000; // mov: $a0 = $t9
hd[241] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[242] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[243] <= 32'b001111_00000_00110_0000000000011110; // li: load 30 in register $a0
hd[244] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[245] <= 32'b001111_00000_01000_0000000000011110; // li: load 30 in register $a2
hd[246] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[247] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[248] <= 32'b011011_11110_00110_0000000000000000; // mov: $a0 = $sp
hd[249] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[250] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[251] <= 32'b001111_00000_00110_0000000000011111; // li: load 31 in register $a0
hd[252] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[253] <= 32'b001111_00000_01000_0000000000011111; // li: load 31 in register $a2
hd[254] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[255] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[256] <= 32'b011011_11111_00110_0000000000000000; // mov: $a0 = $ra
hd[257] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[258] <= 32'b010000_00111_00110_0000000000000000; // sw: mem[$a1 + (0)] = mem[$a0]
hd[259] <= 32'b001111_00000_00110_0000000001000101; // li: load 69 in register $a0
hd[260] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[261] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[262] <= 32'b001100_11110_11110_0000000000000111; // addi: $sp = $sp + (7)
hd[263] <= 32'b010000_11110_00110_1111111111111100; // sw: mem[$sp + (-4)] = mem[$a0]
hd[264] <= 32'b001111_00000_00110_0000000001011001; // li: load 89 in register $a0
hd[265] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[266] <= 32'b100110_00101_01010_0000000000010111; // la: $s0 = mem[$gp + (23)]
hd[267] <= 32'b001110_11110_01011_1111111111111100; // lw: $s1 = mem[$sp] + (-4)
hd[268] <= 32'b000000_01010_01011_10100_00000000000; // add: $t0 = $s0 + $s1
hd[269] <= 32'b001110_10100_10100_0000000000000000; // lw: $t0 = mem[$t0] + (0)
hd[270] <= 32'b010000_11110_10100_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t0]
hd[271] <= 32'b001111_00000_10101_0000000000000000; // li: load 0 in register $t1
hd[272] <= 32'b010000_11110_10101_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t1]
hd[273] <= 32'b001110_00101_01100_0000000000000001; // lw: $s2 = mem[$gp] + (1)
hd[274] <= 32'b000111_01100_01011_10110_00000000000; // mul: $t2 = $s2 * $s1
hd[275] <= 32'b010000_11110_10110_0000000000000000; // sw: mem[$sp + (0)] = mem[$t2]
hd[276] <= 32'b001110_11110_01101_0000000000000000; // lw: $s3 = mem[$sp] + (0)
hd[277] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
hd[278] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[279] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
hd[280] <= 32'b001110_11110_01011_1111111111111101; // lw: $s1 = mem[$sp] + (-3)
hd[281] <= 32'b110000_01010_01011_10111_00000000000; // lt: if($s0 < $s1): $t3 = 1, else $t3 = 0
hd[282] <= 32'b010001_10111_00000_0000000100101010; // bneq: if($t3 == 0) jump to 298
hd[283] <= 32'b001110_11110_01100_0000000000000000; // lw: $s2 = mem[$sp] + (0)
hd[284] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
hd[285] <= 32'b110010_00110_11000_0000000000000000; // lhd: $t4 = hd[$a0]
hd[286] <= 32'b010000_11110_11000_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t4]
hd[287] <= 32'b001110_11110_01101_1111111111111111; // lw: $s3 = mem[$sp] + (-1)
hd[288] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
hd[289] <= 32'b011011_01010_00111_0000000000000000; // mov: $a1 = $s0
hd[290] <= 32'b110111_00111_00110_0000000000000000; // smem_proc: mem[$a0] = $a1
hd[291] <= 32'b001100_01010_11001_0000000000000001; // addi: $t5 = $s0 + (1)
hd[292] <= 32'b010000_11110_11001_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t5]
hd[293] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
hd[294] <= 32'b001100_01100_11010_0000000000000001; // addi: $t6 = $s2 + (1)
hd[295] <= 32'b010000_11110_11010_0000000000000000; // sw: mem[$sp + (0)] = mem[$t6]
hd[296] <= 32'b001110_11110_01100_0000000000000000; // lw: $s2 = mem[$sp] + (0)
hd[297] <= 32'b011010_00000000000000000100010111; // jump to 279 (L1)
hd[298] <= 32'b001110_11110_01010_1111111111111100; // lw: $s0 = mem[$sp] + (-4)
hd[299] <= 32'b001100_01010_11011_0000000000000001; // addi: $t7 = $s0 + (1)
hd[300] <= 32'b010000_11110_11011_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t7]
hd[301] <= 32'b001110_11110_01010_1111111111111100; // lw: $s0 = mem[$sp] + (-4)
hd[302] <= 32'b001110_00101_01011_0000000000000001; // lw: $s1 = mem[$gp] + (1)
hd[303] <= 32'b000111_01010_01011_11100_00000000000; // mul: $t8 = $s0 * $s1
hd[304] <= 32'b010000_11110_11100_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t8]
hd[305] <= 32'b001111_00000_00110_0000000000000001; // li: load 1 in register $a0
hd[306] <= 32'b001110_11110_01100_1111111111111110; // lw: $s2 = mem[$sp] + (-2)
hd[307] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[308] <= 32'b001111_00000_01000_0000000000000001; // li: load 1 in register $a2
hd[309] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[310] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[311] <= 32'b001110_00111_00001_0000000000000000; // lw: $v0 = mem[$a1] + (0)
hd[312] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[313] <= 32'b001111_00000_00110_0000000000000010; // li: load 2 in register $a0
hd[314] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[315] <= 32'b001111_00000_01000_0000000000000010; // li: load 2 in register $a2
hd[316] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[317] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[318] <= 32'b001110_00111_00010_0000000000000000; // lw: $v1 = mem[$a1] + (0)
hd[319] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[320] <= 32'b001111_00000_00110_0000000000000011; // li: load 3 in register $a0
hd[321] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[322] <= 32'b001111_00000_01000_0000000000000011; // li: load 3 in register $a2
hd[323] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[324] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[325] <= 32'b001110_00111_00011_0000000000000000; // lw: $out1 = mem[$a1] + (0)
hd[326] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[327] <= 32'b001111_00000_00110_0000000000000100; // li: load 4 in register $a0
hd[328] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[329] <= 32'b001111_00000_01000_0000000000000100; // li: load 4 in register $a2
hd[330] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[331] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[332] <= 32'b001110_00111_00100_0000000000000000; // lw: $out2 = mem[$a1] + (0)
hd[333] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[334] <= 32'b001111_00000_00110_0000000000000101; // li: load 5 in register $a0
hd[335] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[336] <= 32'b001111_00000_01000_0000000000000101; // li: load 5 in register $a2
hd[337] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[338] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[339] <= 32'b001110_00111_00101_0000000000000000; // lw: $gp = mem[$a1] + (0)
hd[340] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[341] <= 32'b001111_00000_00110_0000000000000110; // li: load 6 in register $a0
hd[342] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[343] <= 32'b001111_00000_01000_0000000000000110; // li: load 6 in register $a2
hd[344] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[345] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[346] <= 32'b001110_00111_00110_0000000000000000; // lw: $a0 = mem[$a1] + (0)
hd[347] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[348] <= 32'b001111_00000_00110_0000000000000111; // li: load 7 in register $a0
hd[349] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[350] <= 32'b001111_00000_01000_0000000000000111; // li: load 7 in register $a2
hd[351] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[352] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[353] <= 32'b001110_00111_00111_0000000000000000; // lw: $a1 = mem[$a1] + (0)
hd[354] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[355] <= 32'b001111_00000_00110_0000000000001000; // li: load 8 in register $a0
hd[356] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[357] <= 32'b001111_00000_01000_0000000000001000; // li: load 8 in register $a2
hd[358] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[359] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[360] <= 32'b001110_00111_01000_0000000000000000; // lw: $a2 = mem[$a1] + (0)
hd[361] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[362] <= 32'b001111_00000_00110_0000000000001001; // li: load 9 in register $a0
hd[363] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[364] <= 32'b001111_00000_01000_0000000000001001; // li: load 9 in register $a2
hd[365] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[366] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[367] <= 32'b001110_00111_01001_0000000000000000; // lw: $a3 = mem[$a1] + (0)
hd[368] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[369] <= 32'b001111_00000_00110_0000000000001010; // li: load 10 in register $a0
hd[370] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[371] <= 32'b001111_00000_01000_0000000000001010; // li: load 10 in register $a2
hd[372] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[373] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[374] <= 32'b001110_00111_01010_0000000000000000; // lw: $s0 = mem[$a1] + (0)
hd[375] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[376] <= 32'b001111_00000_00110_0000000000001011; // li: load 11 in register $a0
hd[377] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[378] <= 32'b001111_00000_01000_0000000000001011; // li: load 11 in register $a2
hd[379] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[380] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[381] <= 32'b001110_00111_01011_0000000000000000; // lw: $s1 = mem[$a1] + (0)
hd[382] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[383] <= 32'b001111_00000_00110_0000000000001100; // li: load 12 in register $a0
hd[384] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[385] <= 32'b001111_00000_01000_0000000000001100; // li: load 12 in register $a2
hd[386] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[387] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[388] <= 32'b001110_00111_01100_0000000000000000; // lw: $s2 = mem[$a1] + (0)
hd[389] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[390] <= 32'b001111_00000_00110_0000000000001101; // li: load 13 in register $a0
hd[391] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[392] <= 32'b001111_00000_01000_0000000000001101; // li: load 13 in register $a2
hd[393] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[394] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[395] <= 32'b001110_00111_01101_0000000000000000; // lw: $s3 = mem[$a1] + (0)
hd[396] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[397] <= 32'b001111_00000_00110_0000000000001110; // li: load 14 in register $a0
hd[398] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[399] <= 32'b001111_00000_01000_0000000000001110; // li: load 14 in register $a2
hd[400] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[401] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[402] <= 32'b001110_00111_01110_0000000000000000; // lw: $s4 = mem[$a1] + (0)
hd[403] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[404] <= 32'b001111_00000_00110_0000000000001111; // li: load 15 in register $a0
hd[405] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[406] <= 32'b001111_00000_01000_0000000000001111; // li: load 15 in register $a2
hd[407] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[408] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[409] <= 32'b001110_00111_01111_0000000000000000; // lw: $s5 = mem[$a1] + (0)
hd[410] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[411] <= 32'b001111_00000_00110_0000000000010000; // li: load 16 in register $a0
hd[412] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[413] <= 32'b001111_00000_01000_0000000000010000; // li: load 16 in register $a2
hd[414] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[415] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[416] <= 32'b001110_00111_10000_0000000000000000; // lw: $s6 = mem[$a1] + (0)
hd[417] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[418] <= 32'b001111_00000_00110_0000000000010001; // li: load 17 in register $a0
hd[419] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[420] <= 32'b001111_00000_01000_0000000000010001; // li: load 17 in register $a2
hd[421] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[422] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[423] <= 32'b001110_00111_10001_0000000000000000; // lw: $s7 = mem[$a1] + (0)
hd[424] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[425] <= 32'b001111_00000_00110_0000000000010010; // li: load 18 in register $a0
hd[426] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[427] <= 32'b001111_00000_01000_0000000000010010; // li: load 18 in register $a2
hd[428] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[429] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[430] <= 32'b001110_00111_10010_0000000000000000; // lw: $s8 = mem[$a1] + (0)
hd[431] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[432] <= 32'b001111_00000_00110_0000000000010011; // li: load 19 in register $a0
hd[433] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[434] <= 32'b001111_00000_01000_0000000000010011; // li: load 19 in register $a2
hd[435] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[436] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[437] <= 32'b001110_00111_10011_0000000000000000; // lw: $s9 = mem[$a1] + (0)
hd[438] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[439] <= 32'b001111_00000_00110_0000000000010100; // li: load 20 in register $a0
hd[440] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[441] <= 32'b001111_00000_01000_0000000000010100; // li: load 20 in register $a2
hd[442] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[443] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[444] <= 32'b001110_00111_10100_0000000000000000; // lw: $t0 = mem[$a1] + (0)
hd[445] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[446] <= 32'b001111_00000_00110_0000000000010101; // li: load 21 in register $a0
hd[447] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[448] <= 32'b001111_00000_01000_0000000000010101; // li: load 21 in register $a2
hd[449] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[450] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[451] <= 32'b001110_00111_10101_0000000000000000; // lw: $t1 = mem[$a1] + (0)
hd[452] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[453] <= 32'b001111_00000_00110_0000000000010110; // li: load 22 in register $a0
hd[454] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[455] <= 32'b001111_00000_01000_0000000000010110; // li: load 22 in register $a2
hd[456] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[457] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[458] <= 32'b001110_00111_10110_0000000000000000; // lw: $t2 = mem[$a1] + (0)
hd[459] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[460] <= 32'b001111_00000_00110_0000000000010111; // li: load 23 in register $a0
hd[461] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[462] <= 32'b001111_00000_01000_0000000000010111; // li: load 23 in register $a2
hd[463] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[464] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[465] <= 32'b001110_00111_10111_0000000000000000; // lw: $t3 = mem[$a1] + (0)
hd[466] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[467] <= 32'b001111_00000_00110_0000000000011000; // li: load 24 in register $a0
hd[468] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[469] <= 32'b001111_00000_01000_0000000000011000; // li: load 24 in register $a2
hd[470] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[471] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[472] <= 32'b001110_00111_11000_0000000000000000; // lw: $t4 = mem[$a1] + (0)
hd[473] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[474] <= 32'b001111_00000_00110_0000000000011001; // li: load 25 in register $a0
hd[475] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[476] <= 32'b001111_00000_01000_0000000000011001; // li: load 25 in register $a2
hd[477] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[478] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[479] <= 32'b001110_00111_11001_0000000000000000; // lw: $t5 = mem[$a1] + (0)
hd[480] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[481] <= 32'b001111_00000_00110_0000000000011010; // li: load 26 in register $a0
hd[482] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[483] <= 32'b001111_00000_01000_0000000000011010; // li: load 26 in register $a2
hd[484] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[485] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[486] <= 32'b001110_00111_11010_0000000000000000; // lw: $t6 = mem[$a1] + (0)
hd[487] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[488] <= 32'b001111_00000_00110_0000000000011011; // li: load 27 in register $a0
hd[489] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[490] <= 32'b001111_00000_01000_0000000000011011; // li: load 27 in register $a2
hd[491] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[492] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[493] <= 32'b001110_00111_11011_0000000000000000; // lw: $t7 = mem[$a1] + (0)
hd[494] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[495] <= 32'b001111_00000_00110_0000000000011100; // li: load 28 in register $a0
hd[496] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[497] <= 32'b001111_00000_01000_0000000000011100; // li: load 28 in register $a2
hd[498] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[499] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[500] <= 32'b001110_00111_11100_0000000000000000; // lw: $t8 = mem[$a1] + (0)
hd[501] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[502] <= 32'b001111_00000_00110_0000000000011101; // li: load 29 in register $a0
hd[503] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[504] <= 32'b001111_00000_01000_0000000000011101; // li: load 29 in register $a2
hd[505] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[506] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[507] <= 32'b001110_00111_11101_0000000000000000; // lw: $t9 = mem[$a1] + (0)
hd[508] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[509] <= 32'b001111_00000_00110_0000000000011110; // li: load 30 in register $a0
hd[510] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[511] <= 32'b001111_00000_01000_0000000000011110; // li: load 30 in register $a2
hd[512] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[513] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[514] <= 32'b001110_00111_11110_0000000000000000; // lw: $sp = mem[$a1] + (0)
hd[515] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[516] <= 32'b001111_00000_00110_0000000000011111; // li: load 31 in register $a0
hd[517] <= 32'b011011_01100_00111_0000000000000000; // mov: $a1 = $s2
hd[518] <= 32'b001111_00000_01000_0000000000011111; // li: load 31 in register $a2
hd[519] <= 32'b000001_00111_01000_00111_00000000000; // sub: $a1 = $a1 - $a2
hd[520] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[521] <= 32'b001110_00111_11111_0000000000000000; // lw: $ra = mem[$a1] + (0)
hd[522] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[523] <= 32'b001111_00000_00110_0000000001100011; // li: load 99 in register $a0
hd[524] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[525] <= 32'b001111_00000_00110_0000000001111011; // li: load 123 in register $a0
hd[526] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[527] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[528] <= 32'b001100_11110_11110_0000000000001010; // addi: $sp = $sp + (10)
hd[529] <= 32'b010000_11110_00110_1111111111111001; // sw: mem[$sp + (-7)] = mem[$a0]
hd[530] <= 32'b001111_00000_10100_0000000000000000; // li: load 0 in register $t0
hd[531] <= 32'b010000_11110_10100_1111111111111011; // sw: mem[$sp + (-5)] = mem[$t0]
hd[532] <= 32'b001111_00000_10101_0000000000000000; // li: load 0 in register $t1
hd[533] <= 32'b010000_11110_10101_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t1]
hd[534] <= 32'b001111_00000_10110_0000000000000000; // li: load 0 in register $t2
hd[535] <= 32'b010000_11110_10110_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t2]
hd[536] <= 32'b001111_00000_00110_0000000000000100; // li: load 4 in register $a0
hd[537] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[538] <= 32'b011100_00000000000000000000000000; // nop
hd[539] <= 32'b100101_00000_10111_0000000000000000; // in $t3
hd[540] <= 32'b010000_00101_10111_0000000000000010; // sw: mem[$gp + (2)] = mem[$t3]
hd[541] <= 32'b001110_11110_01010_1111111111111011; // lw: $s0 = mem[$sp] + (-5)
hd[542] <= 32'b001110_11110_01011_1111111111111001; // lw: $s1 = mem[$sp] + (-7)
hd[543] <= 32'b110000_01010_01011_11000_00000000000; // lt: if($s0 < $s1): $t4 = 1, else $t4 = 0
hd[544] <= 32'b010001_11000_00000_0000001010011000; // bneq: if($t4 == 0) jump to 664
hd[545] <= 32'b001111_00000_00110_0000000000001100; // li: load 12 in register $a0
hd[546] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[547] <= 32'b100110_00101_01100_0000000000000011; // la: $s2 = mem[$gp + (3)]
hd[548] <= 32'b001110_11110_01101_1111111111111100; // lw: $s3 = mem[$sp] + (-4)
hd[549] <= 32'b000000_01100_01101_11001_00000000000; // add: $t5 = $s2 + $s3
hd[550] <= 32'b001110_11001_11001_0000000000000000; // lw: $t5 = mem[$t5] + (0)
hd[551] <= 32'b010000_11110_11001_1111111111111010; // sw: mem[$sp + (-6)] = mem[$t5]
hd[552] <= 32'b001110_11110_01110_1111111111111010; // lw: $s4 = mem[$sp] + (-6)
hd[553] <= 32'b010000_11110_01110_1111111111111101; // sw: mem[$sp + (-3)] = mem[$s4]
hd[554] <= 32'b100110_00101_01111_0000000000101011; // la: $s5 = mem[$gp + (43)]
hd[555] <= 32'b001110_11110_10000_1111111111111101; // lw: $s6 = mem[$sp] + (-3)
hd[556] <= 32'b000000_01111_10000_11010_00000000000; // add: $t6 = $s5 + $s6
hd[557] <= 32'b001110_11010_11010_0000000000000000; // lw: $t6 = mem[$t6] + (0)
hd[558] <= 32'b001111_00000_11011_0000000000000000; // li: load 0 in register $t7
hd[559] <= 32'b011110_11010_11011_11100_00000000000; // eq: if($t6 == $t7): $t8 = 1, else $t8 = 0
hd[560] <= 32'b010001_11100_00000_0000001010001100; // bneq: if($t8 == 0) jump to 652
hd[561] <= 32'b011011_10000_00110_0000000000000000; // mov: $a0 = $s6
hd[562] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[563] <= 32'b100110_00101_10001_0000000000100001; // la: $s7 = mem[$gp + (33)]
hd[564] <= 32'b000000_10001_10000_11101_00000000000; // add: $t9 = $s7 + $s6
hd[565] <= 32'b001110_11101_11101_0000000000000000; // lw: $t9 = mem[$t9] + (0)
hd[566] <= 32'b010000_11110_11101_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t9]
hd[567] <= 32'b001110_11110_10010_1111111111111111; // lw: $s8 = mem[$sp] + (-1)
hd[568] <= 32'b011011_10010_00110_0000000000000000; // mov: $a0 = $s8
hd[569] <= 32'b111110_00000_00110_0000000000000000; // process pc = $a0 
hd[570] <= 32'b011011_10000_00110_0000000000000000; // mov: $a0 = $s6
hd[571] <= 32'b010000_11110_11111_1111111111111000; // sw: mem[$sp + (-8)] = mem[$ra]
hd[572] <= 32'b100001_00000000000000000100000110; // jump and link to 262 (load_proc_context)
hd[573] <= 32'b001101_11110_11110_0000000000000111; // subi: $sp = $sp - (7)
hd[574] <= 32'b001110_11110_11111_1111111111111000; // lw: $ra = mem[$sp] + (-8)
hd[575] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[576] <= 32'b001110_11110_01011_1111111111111101; // lw: $s1 = mem[$sp] + (-3)
hd[577] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
hd[578] <= 32'b011100_00000000000000000000000000; // nop
hd[579] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[580] <= 32'b011011_00110_00110_0000000000000000; // mov: $a0 = $a0
hd[581] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[582] <= 32'b011011_00110_10011_0000000000000000; // mov: $s9 = $a0
hd[583] <= 32'b100111_00000_10011_0000000000000000; // sprc = $s9 
hd[584] <= 32'b011100_00000000000000000000000000; // nop
hd[585] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[586] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[587] <= 32'b011100_00000000000000000000000000; // nop
hd[588] <= 32'b001111_00000_00110_0000000001000110; // li: load 70 in register $a0
hd[589] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[590] <= 32'b011011_00010_01100_0000000000000000; // mov: $s2 = $v1
hd[591] <= 32'b010000_11110_01100_0000000000000000; // sw: mem[$sp + (0)] = mem[$s2]
hd[592] <= 32'b001110_11110_01101_0000000000000000; // lw: $s3 = mem[$sp] + (0)
hd[593] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
hd[594] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[595] <= 32'b111101_00000_00000_0000000000000000; // $v1 = process pc
hd[596] <= 32'b011011_00010_01110_0000000000000000; // mov: $s4 = $v1
hd[597] <= 32'b100110_00101_01111_0000000000100001; // la: $s5 = mem[$gp + (33)]
hd[598] <= 32'b000000_01111_01011_10100_00000000000; // add: $t0 = $s5 + $s1
hd[599] <= 32'b010000_10100_01110_0000000000000000; // sw: mem[$t0 + (0)] = mem[$s4]
hd[600] <= 32'b001111_00000_10101_0000000000000001; // li: load 1 in register $t1
hd[601] <= 32'b011110_01101_10101_10110_00000000000; // eq: if($s3 == $t1): $t2 = 1, else $t2 = 0
hd[602] <= 32'b010001_10110_00000_0000001001100111; // bneq: if($t2 == 0) jump to 615
hd[603] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
hd[604] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[605] <= 32'b011100_00000000000000000000000000; // nop
hd[606] <= 32'b100101_00000_10111_0000000000000000; // in $t3
hd[607] <= 32'b010000_11110_10111_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t3]
hd[608] <= 32'b001110_11110_10000_1111111111111110; // lw: $s6 = mem[$sp] + (-2)
hd[609] <= 32'b011011_10000_00110_0000000000000000; // mov: $a0 = $s6
hd[610] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[611] <= 32'b011011_10000_00110_0000000000000000; // mov: $a0 = $s6
hd[612] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[613] <= 32'b011011_00110_00010_0000000000000000; // mov: $v1 = $a0
hd[614] <= 32'b111000_00000_00000_0000000000000000; // chrt
hd[615] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[616] <= 32'b001111_00000_11000_0000000000000010; // li: load 2 in register $t4
hd[617] <= 32'b011110_01010_11000_11001_00000000000; // eq: if($s0 == $t4): $t5 = 1, else $t5 = 0
hd[618] <= 32'b010001_11001_00000_0000001001110100; // bneq: if($t5 == 0) jump to 628
hd[619] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[620] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[621] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[622] <= 32'b011011_00010_01011_0000000000000000; // mov: $s1 = $v1
hd[623] <= 32'b111001_00000_00000_0000000000000000; // chrd
hd[624] <= 32'b010000_11110_01011_1111111111111110; // sw: mem[$sp + (-2)] = mem[$s1]
hd[625] <= 32'b001110_11110_01100_1111111111111110; // lw: $s2 = mem[$sp] + (-2)
hd[626] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
hd[627] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[628] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[629] <= 32'b001111_00000_11010_0000000000000011; // li: load 3 in register $t6
hd[630] <= 32'b011110_01010_11010_11011_00000000000; // eq: if($s0 == $t6): $t7 = 1, else $t7 = 0
hd[631] <= 32'b010001_11011_00000_0000001010000101; // bneq: if($t7 == 0) jump to 645
hd[632] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[633] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[634] <= 32'b001110_11110_01011_1111111111111101; // lw: $s1 = mem[$sp] + (-3)
hd[635] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
hd[636] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[637] <= 32'b100110_00101_01100_0000000000101011; // la: $s2 = mem[$gp + (43)]
hd[638] <= 32'b000000_01100_01011_11100_00000000000; // add: $t8 = $s2 + $s1
hd[639] <= 32'b001111_00000_11101_0000000000000001; // li: load 1 in register $t9
hd[640] <= 32'b010000_11100_11101_0000000000000000; // sw: mem[$t8 + (0)] = mem[$t9]
hd[641] <= 32'b001110_11110_01101_1111111111111011; // lw: $s3 = mem[$sp] + (-5)
hd[642] <= 32'b001100_01101_10100_0000000000000001; // addi: $t0 = $s3 + (1)
hd[643] <= 32'b010000_11110_10100_1111111111111011; // sw: mem[$sp + (-5)] = mem[$t0]
hd[644] <= 32'b001110_11110_01101_1111111111111011; // lw: $s3 = mem[$sp] + (-5)
hd[645] <= 32'b001110_11110_01010_1111111111111101; // lw: $s0 = mem[$sp] + (-3)
hd[646] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[647] <= 32'b010000_11110_11111_1111111111111000; // sw: mem[$sp + (-8)] = mem[$ra]
hd[648] <= 32'b100001_00000000000000000000000001; // jump and link to 1 (store_proc_context)
hd[649] <= 32'b001101_11110_11110_0000000000000100; // subi: $sp = $sp - (4)
hd[650] <= 32'b001110_11110_11111_1111111111111000; // lw: $ra = mem[$sp] + (-8)
hd[651] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[652] <= 32'b001110_11110_01010_1111111111111001; // lw: $s0 = mem[$sp] + (-7)
hd[653] <= 32'b001101_01010_10101_0000000000000001; // subi: $t1 = $s0 - (1)
hd[654] <= 32'b001110_11110_01011_1111111111111100; // lw: $s1 = mem[$sp] + (-4)
hd[655] <= 32'b110000_01011_10101_10110_00000000000; // lt: if($s1 < $t1): $t2 = 1, else $t2 = 0
hd[656] <= 32'b010001_10110_00000_0000001010010101; // bneq: if($t2 == 0) jump to 661
hd[657] <= 32'b001100_01011_10111_0000000000000001; // addi: $t3 = $s1 + (1)
hd[658] <= 32'b010000_11110_10111_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t3]
hd[659] <= 32'b001110_11110_01011_1111111111111100; // lw: $s1 = mem[$sp] + (-4)
hd[660] <= 32'b011010_00000000000000001010010111; // jump to 663 (L9)
hd[661] <= 32'b001111_00000_11000_0000000000000000; // li: load 0 in register $t4
hd[662] <= 32'b010000_11110_11000_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t4]
hd[663] <= 32'b011010_00000000000000001000011101; // jump to 541 (L3)
hd[664] <= 32'b001111_00000_00110_0000000000000101; // li: load 5 in register $a0
hd[665] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[666] <= 32'b011100_00000000000000000000000000; // nop
hd[667] <= 32'b100101_00000_11001_0000000000000000; // in $t5
hd[668] <= 32'b010000_00101_11001_0000000000000010; // sw: mem[$gp + (2)] = mem[$t5]
hd[669] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[670] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
hd[671] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[672] <= 32'b001111_00000_10100_0000000000001010; // li: load 10 in register $t0
hd[673] <= 32'b110000_01010_10100_10101_00000000000; // lt: if($s0 < $t0): $t1 = 1, else $t1 = 0
hd[674] <= 32'b010001_10101_00000_0000001010101011; // bneq: if($t1 == 0) jump to 683
hd[675] <= 32'b100110_00101_01011_0000000000000011; // la: $s1 = mem[$gp + (3)]
hd[676] <= 32'b000000_01011_01010_10110_00000000000; // add: $t2 = $s1 + $s0
hd[677] <= 32'b001111_00000_10111_0000000000000000; // li: load 0 in register $t3
hd[678] <= 32'b010000_10110_10111_0000000000000000; // sw: mem[$t2 + (0)] = mem[$t3]
hd[679] <= 32'b001100_01010_11000_0000000000000001; // addi: $t4 = $s0 + (1)
hd[680] <= 32'b010000_11110_11000_0000000000000000; // sw: mem[$sp + (0)] = mem[$t4]
hd[681] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[682] <= 32'b011010_00000000000000001010011111; // jump to 671 (L11)
hd[683] <= 32'b001111_00000_00110_0000000001010111; // li: load 87 in register $a0
hd[684] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[685] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[686] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
hd[687] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[688] <= 32'b001111_00000_10100_0000000000001010; // li: load 10 in register $t0
hd[689] <= 32'b110000_01010_10100_10101_00000000000; // lt: if($s0 < $t0): $t1 = 1, else $t1 = 0
hd[690] <= 32'b010001_10101_00000_0000001010111011; // bneq: if($t1 == 0) jump to 699
hd[691] <= 32'b100110_00101_01011_0000000000100001; // la: $s1 = mem[$gp + (33)]
hd[692] <= 32'b000000_01011_01010_10110_00000000000; // add: $t2 = $s1 + $s0
hd[693] <= 32'b001111_00000_10111_0000000000000000; // li: load 0 in register $t3
hd[694] <= 32'b010000_10110_10111_0000000000000000; // sw: mem[$t2 + (0)] = mem[$t3]
hd[695] <= 32'b001100_01010_11000_0000000000000001; // addi: $t4 = $s0 + (1)
hd[696] <= 32'b010000_11110_11000_0000000000000000; // sw: mem[$sp + (0)] = mem[$t4]
hd[697] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[698] <= 32'b011010_00000000000000001010101111; // jump to 687 (L13)
hd[699] <= 32'b001111_00000_00110_0000000000101111; // li: load 47 in register $a0
hd[700] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[701] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[702] <= 32'b001100_11110_11110_0000000000000101; // addi: $sp = $sp + (5)
hd[703] <= 32'b001111_00000_00110_0000000000000010; // li: load 2 in register $a0
hd[704] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[705] <= 32'b011100_00000000000000000000000000; // nop
hd[706] <= 32'b100101_00000_10100_0000000000000000; // in $t0
hd[707] <= 32'b010000_11110_10100_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t0]
hd[708] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
hd[709] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[710] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[711] <= 32'b001111_00000_10101_0000000000000000; // li: load 0 in register $t1
hd[712] <= 32'b010000_11110_10101_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t1]
hd[713] <= 32'b001111_00000_00110_0000000000000011; // li: load 3 in register $a0
hd[714] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[715] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[716] <= 32'b001110_11110_01011_1111111111111110; // lw: $s1 = mem[$sp] + (-2)
hd[717] <= 32'b110000_01010_01011_10110_00000000000; // lt: if($s0 < $s1): $t2 = 1, else $t2 = 0
hd[718] <= 32'b010001_10110_00000_0000001011100000; // bneq: if($t2 == 0) jump to 736
hd[719] <= 32'b011100_00000000000000000000000000; // nop
hd[720] <= 32'b100101_00000_10111_0000000000000000; // in $t3
hd[721] <= 32'b010000_11110_10111_0000000000000000; // sw: mem[$sp + (0)] = mem[$t3]
hd[722] <= 32'b001110_11110_01100_0000000000000000; // lw: $s2 = mem[$sp] + (0)
hd[723] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
hd[724] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[725] <= 32'b100110_00101_01101_0000000000000011; // la: $s3 = mem[$gp + (3)]
hd[726] <= 32'b000000_01101_01010_11000_00000000000; // add: $t4 = $s3 + $s0
hd[727] <= 32'b010000_11000_01100_0000000000000000; // sw: mem[$t4 + (0)] = mem[$s2]
hd[728] <= 32'b100110_00101_01110_0000000000101011; // la: $s4 = mem[$gp + (43)]
hd[729] <= 32'b000000_01110_01010_11001_00000000000; // add: $t5 = $s4 + $s0
hd[730] <= 32'b001111_00000_11010_0000000000000000; // li: load 0 in register $t6
hd[731] <= 32'b010000_11001_11010_0000000000000000; // sw: mem[$t5 + (0)] = mem[$t6]
hd[732] <= 32'b001100_01010_11011_0000000000000001; // addi: $t7 = $s0 + (1)
hd[733] <= 32'b010000_11110_11011_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t7]
hd[734] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[735] <= 32'b011010_00000000000000001011001011; // jump to 715 (L15)
hd[736] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
hd[737] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[738] <= 32'b010000_11110_11111_1111111111111101; // sw: mem[$sp + (-3)] = mem[$ra]
hd[739] <= 32'b100001_00000000000000001000010000; // jump and link to 528 (circular_queue)
hd[740] <= 32'b001101_11110_11110_0000000000001010; // subi: $sp = $sp - (10)
hd[741] <= 32'b001110_11110_11111_1111111111111101; // lw: $ra = mem[$sp] + (-3)
hd[742] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[743] <= 32'b010000_11110_11111_1111111111111101; // sw: mem[$sp + (-3)] = mem[$ra]
hd[744] <= 32'b100001_00000000000000001010011110; // jump and link to 670 (reset_queue)
hd[745] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
hd[746] <= 32'b001110_11110_11111_1111111111111101; // lw: $ra = mem[$sp] + (-3)
hd[747] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[748] <= 32'b010000_11110_11111_1111111111111101; // sw: mem[$sp + (-3)] = mem[$ra]
hd[749] <= 32'b100001_00000000000000001010101110; // jump and link to 686 (reset_pcs)
hd[750] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
hd[751] <= 32'b001110_11110_11111_1111111111111101; // lw: $ra = mem[$sp] + (-3)
hd[752] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[753] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[754] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
hd[755] <= 32'b001111_00000_00110_0000000000000001; // li: load 1 in register $a0
hd[756] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[757] <= 32'b011100_00000000000000000000000000; // nop
hd[758] <= 32'b100101_00000_10100_0000000000000000; // in $t0
hd[759] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
hd[760] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[761] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
hd[762] <= 32'b111111_00000_00110_0000000000000000; // out $a0
hd[763] <= 32'b001111_00000_10101_0000000000000001; // li: load 1 in register $t1
hd[764] <= 32'b011110_01010_10101_10110_00000000000; // eq: if($s0 == $t1): $t2 = 1, else $t2 = 0
hd[765] <= 32'b010001_10110_00000_0000001100000011; // bneq: if($t2 == 0) jump to 771
hd[766] <= 32'b010000_11110_11111_1111111111111111; // sw: mem[$sp + (-1)] = mem[$ra]
hd[767] <= 32'b100001_00000000000000001010111110; // jump and link to 702 (process_handling)
hd[768] <= 32'b001101_11110_11110_0000000000000101; // subi: $sp = $sp - (5)
hd[769] <= 32'b001110_11110_11111_1111111111111111; // lw: $ra = mem[$sp] + (-1)
hd[770] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[771] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[772] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
hd[773] <= 32'b001111_00000_10100_0000000000000000; // li: load 0 in register $t0
hd[774] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
hd[775] <= 32'b001111_00000_10101_0000000000001010; // li: load 10 in register $t1
hd[776] <= 32'b010000_00101_10101_0000000000000000; // sw: mem[$gp + (0)] = mem[$t1]
hd[777] <= 32'b001111_00000_10110_0000010000000000; // li: load 1024 in register $t2
hd[778] <= 32'b010000_00101_10110_0000000000000001; // sw: mem[$gp + (1)] = mem[$t2]
hd[779] <= 32'b100110_00101_01010_0000000000010111; // la: $s0 = mem[$gp + (23)]
hd[780] <= 32'b001111_00000_10111_0000000000110010; // li: load 50 in register $t3
hd[781] <= 32'b010000_01010_10111_0000000000000001; // sw: mem[$s0 + (1)] = mem[$t3]
hd[782] <= 32'b001111_00000_11000_0000000000110010; // li: load 50 in register $t4
hd[783] <= 32'b010000_01010_11000_0000000000000010; // sw: mem[$s0 + (2)] = mem[$t4]
hd[784] <= 32'b001111_00000_11001_0000000000110010; // li: load 50 in register $t5
hd[785] <= 32'b010000_01010_11001_0000000000000011; // sw: mem[$s0 + (3)] = mem[$t5]
hd[786] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[787] <= 32'b001111_00000_11010_0000000000001010; // li: load 10 in register $t6
hd[788] <= 32'b110000_01010_11010_11011_00000000000; // lt: if($s0 < $t6): $t7 = 1, else $t7 = 0
hd[789] <= 32'b010001_11011_00000_0000001100101001; // bneq: if($t7 == 0) jump to 809
hd[790] <= 32'b100110_00101_01011_0000000000000011; // la: $s1 = mem[$gp + (3)]
hd[791] <= 32'b000000_01011_01010_11100_00000000000; // add: $t8 = $s1 + $s0
hd[792] <= 32'b001111_00000_11101_0000000000000000; // li: load 0 in register $t9
hd[793] <= 32'b010000_11100_11101_0000000000000000; // sw: mem[$t8 + (0)] = mem[$t9]
hd[794] <= 32'b100110_00101_01100_0000000000101011; // la: $s2 = mem[$gp + (43)]
hd[795] <= 32'b000000_01100_01010_10100_00000000000; // add: $t0 = $s2 + $s0
hd[796] <= 32'b001111_00000_10101_0000000000000000; // li: load 0 in register $t1
hd[797] <= 32'b010000_10100_10101_0000000000000000; // sw: mem[$t0 + (0)] = mem[$t1]
hd[798] <= 32'b100110_00101_01101_0000000000100001; // la: $s3 = mem[$gp + (33)]
hd[799] <= 32'b000000_01101_01010_10110_00000000000; // add: $t2 = $s3 + $s0
hd[800] <= 32'b001111_00000_10111_0000000000000000; // li: load 0 in register $t3
hd[801] <= 32'b010000_10110_10111_0000000000000000; // sw: mem[$t2 + (0)] = mem[$t3]
hd[802] <= 32'b100110_00101_01110_0000000000001101; // la: $s4 = mem[$gp + (13)]
hd[803] <= 32'b000000_01110_01010_11000_00000000000; // add: $t4 = $s4 + $s0
hd[804] <= 32'b010000_11000_01010_0000000000000000; // sw: mem[$t4 + (0)] = mem[$s0]
hd[805] <= 32'b001100_01010_11001_0000000000000001; // addi: $t5 = $s0 + (1)
hd[806] <= 32'b010000_11110_11001_0000000000000000; // sw: mem[$sp + (0)] = mem[$t5]
hd[807] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[808] <= 32'b011010_00000000000000001100010010; // jump to 786 (L18)
hd[809] <= 32'b011001_11111_00000_00000_00000000000; // jr: jump to register $ra
hd[810] <= 32'b001100_00101_11110_0000000000000001; // addi: $sp = $gp + (1)
hd[811] <= 32'b001100_11110_11110_0000000000110110; // addi: $sp = $sp + (54)
hd[812] <= 32'b010000_11110_11111_0000000000000000; // sw: mem[$sp + (0)] = mem[$ra]
hd[813] <= 32'b100001_00000000000000001100000100; // jump and link to 772 (init_os)
hd[814] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
hd[815] <= 32'b001110_11110_11111_0000000000000000; // lw: $ra = mem[$sp] + (0)
hd[816] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[817] <= 32'b001111_00000_00110_0000000000000000; // li: load 0 in register $a0
hd[818] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
hd[819] <= 32'b011100_00000000000000000000000000; // nop
hd[820] <= 32'b100101_00000_10100_0000000000000000; // in $t0
hd[821] <= 32'b010000_00101_10100_0000000000000010; // sw: mem[$gp + (2)] = mem[$t0]
hd[822] <= 32'b001111_00000_10101_0000000000000001; // li: load 1 in register $t1
hd[823] <= 32'b001111_00000_10110_0000000000000010; // li: load 2 in register $t2
hd[824] <= 32'b110000_10101_10110_10111_00000000000; // lt: if($t1 < $t2): $t3 = 1, else $t3 = 0
hd[825] <= 32'b010001_10111_00000_0000001101000000; // bneq: if($t3 == 0) jump to 832
hd[826] <= 32'b010000_11110_11111_0000000000000000; // sw: mem[$sp + (0)] = mem[$ra]
hd[827] <= 32'b100001_00000000000000001011110010; // jump and link to 754 (bash)
hd[828] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
hd[829] <= 32'b001110_11110_11111_0000000000000000; // lw: $ra = mem[$sp] + (0)
hd[830] <= 32'b011011_00001_01010_0000000000000000; // mov: $s0 = $v0
hd[831] <= 32'b011010_00000000000000001100110110; // jump to 822 (L20)
hd[832] <= 32'b001101_11110_11110_0000000000000001; // subi: $sp = $sp - (1)
hd[833] <= 32'b011101_00000000000000000000000000; // hlt










//processes
//prog1
hd[1024] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
hd[1025] <= 32'b001100_11110_11110_0000000000000100; // addi: $sp = $sp + (4)
hd[1026] <= 32'b011100_00000000000000000000000000; // nop
hd[1027] <= 32'b111010_00000000000000000000000000; // sysin
hd[1028] <= 32'b011100_00000000000000000000000000; // nop
hd[1029] <= 32'b011100_00000000000000000000000000; // nop
hd[1030] <= 32'b010000_11110_00010_1111111111111110; // sw: mem[$sp + (-2)] = mem[$v1]
hd[1031] <= 32'b001110_11110_01010_1111111111111110; // lw: $s0 = mem[$sp] + (-2)
hd[1032] <= 32'b001100_01010_10101_0000000000001101; // addi: $t1 = $s0 + (13)
hd[1033] <= 32'b010000_11110_10101_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t1]
hd[1034] <= 32'b001110_11110_01011_1111111111111111; // lw: $s1 = mem[$sp] + (-1)
hd[1035] <= 32'b011011_01011_00010_0000000000000000; // mov: $v1 = $s1
hd[1036] <= 32'b011100_00000000000000000000000000; // nop
hd[1037] <= 32'b111011_00000000000000000000000000; // sysout
hd[1038] <= 32'b011100_00000000000000000000000000; // nop
hd[1039] <= 32'b001101_11110_11110_0000000000000100; // subi: $sp = $sp - (4)
hd[1040] <= 32'b111100_00000000000000000000000000; // sysend
hd[1041] <= 32'b011100_00000000000000000000000000; // nop

//prog2
hd[2048] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
hd[2049] <= 32'b001100_11110_11110_0000000000000111; // addi: $sp = $sp + (7)
hd[2050] <= 32'b011100_00000000000000000000000000; // nop
hd[2051] <= 32'b111010_00000000000000000000000000; // sysin
hd[2052] <= 32'b011100_00000000000000000000000000; // nop
hd[2053] <= 32'b011100_00000000000000000000000000; // nop
hd[2054] <= 32'b010000_11110_00010_1111111111111011; // sw: mem[$sp + (-5)] = mem[$v1]
hd[2055] <= 32'b001110_11110_01010_1111111111111011; // lw: $s0 = mem[$sp] + (-5)
hd[2056] <= 32'b001100_01010_10101_0000000000000001; // addi: $t1 = $s0 + (1)
hd[2057] <= 32'b010000_11110_10101_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t1]
hd[2058] <= 32'b001110_11110_01011_1111111111111100; // lw: $s1 = mem[$sp] + (-4)
hd[2059] <= 32'b001100_01011_10110_0000000000000001; // addi: $t2 = $s1 + (1)
hd[2060] <= 32'b010000_11110_10110_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t2]
hd[2061] <= 32'b001110_11110_01100_1111111111111101; // lw: $s2 = mem[$sp] + (-3)
hd[2062] <= 32'b011011_01100_00010_0000000000000000; // mov: $v1 = $s2
hd[2063] <= 32'b011100_00000000000000000000000000; // nop
hd[2064] <= 32'b111011_00000000000000000000000000; // sysout
hd[2065] <= 32'b011100_00000000000000000000000000; // nop
hd[2066] <= 32'b001101_11110_11110_0000000000000111; // subi: $sp = $sp - (7)
hd[2067] <= 32'b111100_00000000000000000000000000; // sysend
hd[2068] <= 32'b011100_00000000000000000000000000; // nop

//prog3

hd[3072] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
hd[3073] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
hd[3074] <= 32'b001111_00000_10100_0000000000000001; // li: load 1 in register $t0
hd[3075] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
hd[3076] <= 32'b011100_00000000000000000000000000; // nop
hd[3077] <= 32'b111010_00000000000000000000000000; // sysin
hd[3078] <= 32'b011100_00000000000000000000000000; // nop
hd[3079] <= 32'b011100_00000000000000000000000000; // nop
hd[3080] <= 32'b010000_11110_00010_1111111111111111; // sw: mem[$sp + (-1)] = mem[$v1]
hd[3081] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[3082] <= 32'b001111_00000_10110_0000000000000000; // li: load 0 in register $t2
hd[3083] <= 32'b100000_01010_10110_10111_00000000000; // gt: if($s0 > $t2): $t3 = 1, else $t3 = 0
hd[3084] <= 32'b010001_10111_00000_0000000000010011; // bneq: if($t3 == 0) jump to 19
hd[3085] <= 32'b000111_01010_01010_11000_00000000000; // mul: $t4 = $s0 * $s0
hd[3086] <= 32'b010000_11110_11000_0000000000000000; // sw: mem[$sp + (0)] = mem[$t4]
hd[3087] <= 32'b001101_01010_11001_0000000000000001; // subi: $t5 = $s0 - (1)
hd[3088] <= 32'b010000_11110_11001_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t5]
hd[3089] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
hd[3090] <= 32'b011010_00000000000000000000001001; // jump to 9 (L1)
hd[3091] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
hd[3092] <= 32'b011011_01010_00010_0000000000000000; // mov: $v1 = $s0
hd[3093] <= 32'b011100_00000000000000000000000000; // nop
hd[3094] <= 32'b111011_00000000000000000000000000; // sysout
hd[3095] <= 32'b011100_00000000000000000000000000; // nop
hd[3096] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
hd[3097] <= 32'b111100_00000000000000000000000000; // sysend
hd[3098] <= 32'b011100_00000000000000000000000000; // nop



	end
	
	always @ ( posedge clk )
	begin
		if( write_flag )
			hd[address] <= input_data; //write to disk
	end
	
	always @ ( posedge clk_auto )
	begin
		hd_output <= hd[address];
	end

endmodule 

	