module BIOS(address, biosOut, clk_auto);

	input [31:0]address;
	input clk_auto;
	output reg [31:0]biosOut;
	
	reg [31:0] bios[63:0];
	initial
		begin				
bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000011; // addi: $sp = $sp + (3)
bios[2] <= 32'b001111_00000_10100_0000000000000000; // li: load 0 in register $t0
bios[3] <= 32'b010000_11110_10100_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t0]
bios[4] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[5] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[6] <= 32'b110010_00110_10101_0000000000000000; // lhd: $t1 = hd[$a0]
bios[7] <= 32'b010000_11110_10101_0000000000000000; // sw: mem[$sp + (0)] = mem[$t1]
bios[8] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[9] <= 32'b001111_00000_10110_0000000100000000; // li: load 256 in register $t2
bios[10] <= 32'b100010_01010_10110_10111_00000000000; // neq: if($s0 != $t2): $t3 = 1, else $t3 = 0
bios[11] <= 32'b010001_10111_00000_0000000000011000; // bneq: if($t3 == 0) jump to 24
bios[12] <= 32'b001110_11110_01011_0000000000000000; // lw: $s1 = mem[$sp] + (0)
bios[13] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
bios[14] <= 32'b011011_01010_00111_0000000000000000; // mov: $a1 = $s0
bios[15] <= 32'b110101_00111_00110_0000000000000000; // smem: mem[$a0] = $a1
bios[16] <= 32'b001100_01010_11000_0000000000000001; // addi: $t4 = $s0 + (1)
bios[17] <= 32'b010000_11110_11000_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t4]
bios[18] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[19] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[20] <= 32'b110010_00110_11001_0000000000000000; // lhd: $t5 = hd[$a0]
bios[21] <= 32'b010000_11110_11001_0000000000000000; // sw: mem[$sp + (0)] = mem[$t5]
bios[22] <= 32'b001110_11110_01011_0000000000000000; // lw: $s1 = mem[$sp] + (0)
bios[23] <= 32'b011010_00000000000000000000001000; // jump to 8 (L1)
bios[24] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
bios[25] <= 32'b011011_01010_00110_0000000000000000; // mov: $a0 = $s0
bios[26] <= 32'b001110_11110_01011_1111111111111111; // lw: $s1 = mem[$sp] + (-1)
bios[27] <= 32'b011011_01011_00111_0000000000000000; // mov: $a1 = $s1
bios[28] <= 32'b110101_00111_00110_0000000000000000; // smem: mem[$a0] = $a1
bios[29] <= 32'b001111_00000_00110_0000000000001000; // li: load 8 in register $a0
bios[30] <= 32'b110110_00000_00110_0000000000000000; // lcd ($a0)
bios[31] <= 32'b011011_01011_00110_0000000000000000; // mov: $a0 = $s1
bios[32] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[33] <= 32'b001111_00000_00110_0000000001100011; // li: load 99 in register $a0
bios[34] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[35] <= 32'b001101_11110_11110_0000000000000011; // subi: $sp = $sp - (3)
bios[36] <= 32'b011101_00000000000000000000000000; // hlt



		end
	
	always @(posedge clk_auto)
		begin
			biosOut <= bios[address];
		end

	
endmodule

