module BIOS(address, biosOut, clk_auto);

	input [31:0]address;
	input clk_auto;
	output reg [31:0]biosOut;
	
	reg [31:0] bios[63:0];
	initial
		begin
		
		
bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000110; // addi: $sp = $sp + (6)
bios[2] <= 32'b001111_00000_10100_0000000011111010; // li: load 250 in register $t0
bios[3] <= 32'b010000_11110_10100_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t0]
bios[4] <= 32'b001111_00000_10101_0000001111101000; // li: load 1000 in register $t1
bios[5] <= 32'b010000_11110_10101_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t1]
bios[6] <= 32'b001110_11110_01010_1111111111111111; // lw: $s0 = mem[$sp] + (-1)
bios[7] <= 32'b001110_11110_01011_1111111111111110; // lw: $s1 = mem[$sp] + (-2)
bios[8] <= 32'b000111_01010_01011_10110_00000000000; // mul: $t2 = $s0 * $s1
bios[9] <= 32'b010000_11110_10110_1111111111111100; // sw: mem[$sp + (-4)] = mem[$t2]
bios[10] <= 32'b001110_11110_01100_1111111111111100; // lw: $s2 = mem[$sp] + (-4)
bios[11] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
bios[12] <= 32'b101101_00000_00110_0000000000000000; // baud $a0
bios[13] <= 32'b011100_00000000000000000000000000; // nop
bios[14] <= 32'b011100_00000000000000000000000000; // nop
bios[15] <= 32'b011100_00000000000000000000000000; // nop
bios[16] <= 32'b011100_00000000000000000000000000; // nop
bios[17] <= 32'b011100_00000000000000000000000000; // nop
bios[18] <= 32'b011100_00000000000000000000000000; // nop
bios[19] <= 32'b011100_00000000000000000000000000; // nop
bios[20] <= 32'b011100_00000000000000000000000000; // nop
bios[21] <= 32'b011100_00000000000000000000000000; // nop
bios[22] <= 32'b011100_00000000000000000000000000; // nop
bios[23] <= 32'b011100_00000000000000000000000000; // nop
bios[24] <= 32'b011100_00000000000000000000000000; // nop
bios[25] <= 32'b011100_00000000000000000000000000; // nop
bios[26] <= 32'b011100_00000000000000000000000000; // nop
bios[27] <= 32'b011100_00000000000000000000000000; // nop
bios[28] <= 32'b011100_00000000000000000000000000; // nop
bios[29] <= 32'b101111_00000_10111_0000000000000000; // rcv $t3
bios[30] <= 32'b010000_11110_10111_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t3]
bios[31] <= 32'b001110_11110_01101_1111111111111101; // lw: $s3 = mem[$sp] + (-3)
bios[32] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
bios[33] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[34] <= 32'b001100_01101_11000_0000000000001100; // addi: $t4 = $s3 + (12)
bios[35] <= 32'b010000_11110_11000_0000000000000000; // sw: mem[$sp + (0)] = mem[$t4]
bios[36] <= 32'b001110_11110_01110_0000000000000000; // lw: $s4 = mem[$sp] + (0)
bios[37] <= 32'b011011_01110_00110_0000000000000000; // mov: $a0 = $s4
bios[38] <= 32'b011100_00000000000000000000000000; // nop
bios[39] <= 32'b011100_00000000000000000000000000; // nop
bios[40] <= 32'b011100_00000000000000000000000000; // nop
bios[41] <= 32'b011100_00000000000000000000000000; // nop
bios[42] <= 32'b011100_00000000000000000000000000; // nop
bios[43] <= 32'b011100_00000000000000000000000000; // nop
bios[44] <= 32'b101110_00000_00110_0000000000000000; // snd $a0
bios[45] <= 32'b001101_11110_11110_0000000000000110; // subi: $sp = $sp - (6)
bios[46] <= 32'b011101_00000000000000000000000000; // hlt


		
/*bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000101; // addi: $sp = $sp + (5)
bios[2] <= 32'b001111_00000_10100_0000000011111010; // li: load 250 in register $t0
bios[3] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
bios[4] <= 32'b001111_00000_10101_0000001111101000; // li: load 1000 in register $t1
bios[5] <= 32'b010000_11110_10101_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t1]
bios[6] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
bios[7] <= 32'b001110_11110_01011_1111111111111111; // lw: $s1 = mem[$sp] + (-1)
bios[8] <= 32'b000111_01010_01011_10110_00000000000; // mul: $t2 = $s0 * $s1
bios[9] <= 32'b010000_11110_10110_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t2]
bios[10] <= 32'b001110_11110_01100_1111111111111101; // lw: $s2 = mem[$sp] + (-3)
bios[11] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
bios[12] <= 32'b101101_00000_00110_0000000000000000; // baud $a0
bios[13] <= 32'b001111_00000_00110_0000000001011000; // li: load 88 in register $a0
bios[14] <= 32'b011100_00000000000000000000000000; // nop
bios[15] <= 32'b011100_00000000000000000000000000; // nop
bios[16] <= 32'b011100_00000000000000000000000000; // nop
bios[17] <= 32'b011100_00000000000000000000000000; // nop
bios[18] <= 32'b011100_00000000000000000000000000; // nop
bios[19] <= 32'b011100_00000000000000000000000000; // nop
bios[20] <= 32'b101110_00000_00110_0000000000000000; // snd $a0
bios[21] <= 32'b001101_11110_11110_0000000000000101; // subi: $sp = $sp - (5)
bios[22] <= 32'b011101_00000000000000000000000000; // hlt*/
		
/*bios[0] <= 32'b011010_00000000000000000000000001; // jump to 1 (main)
bios[1] <= 32'b001100_11110_11110_0000000000000101; // addi: $sp = $sp + (5)
bios[2] <= 32'b001111_00000_10100_0000000011111010; // li: load 250 in register $t0
bios[3] <= 32'b010000_11110_10100_0000000000000000; // sw: mem[$sp + (0)] = mem[$t0]
bios[4] <= 32'b001111_00000_10101_0000001111101000; // li: load 1000 in register $t1
bios[5] <= 32'b010000_11110_10101_1111111111111111; // sw: mem[$sp + (-1)] = mem[$t1]
bios[6] <= 32'b001110_11110_01010_0000000000000000; // lw: $s0 = mem[$sp] + (0)
bios[7] <= 32'b001110_11110_01011_1111111111111111; // lw: $s1 = mem[$sp] + (-1)
bios[8] <= 32'b000111_01010_01011_10110_00000000000; // mul: $t2 = $s0 * $s1
bios[9] <= 32'b010000_11110_10110_1111111111111101; // sw: mem[$sp + (-3)] = mem[$t2]
bios[10] <= 32'b001110_11110_01100_1111111111111101; // lw: $s2 = mem[$sp] + (-3)
bios[11] <= 32'b011011_01100_00110_0000000000000000; // mov: $a0 = $s2
bios[12] <= 32'b101101_00000_00110_0000000000000000; // baud $a0
bios[13] <= 32'b011100_00000000000000000000000000; // nop
bios[14] <= 32'b011100_00000000000000000000000000; // nop
bios[15] <= 32'b011100_00000000000000000000000000; // nop
bios[16] <= 32'b011100_00000000000000000000000000; // nop
bios[17] <= 32'b011100_00000000000000000000000000; // nop
bios[18] <= 32'b011100_00000000000000000000000000; // nop
bios[19] <= 32'b011100_00000000000000000000000000; // nop
bios[20] <= 32'b011100_00000000000000000000000000; // nop
bios[21] <= 32'b011100_00000000000000000000000000; // nop
bios[22] <= 32'b011100_00000000000000000000000000; // nop
bios[23] <= 32'b011100_00000000000000000000000000; // nop
bios[24] <= 32'b011100_00000000000000000000000000; // nop
bios[25] <= 32'b011100_00000000000000000000000000; // nop
bios[26] <= 32'b011100_00000000000000000000000000; // nop
bios[27] <= 32'b011100_00000000000000000000000000; // nop
bios[28] <= 32'b011100_00000000000000000000000000; // nop
bios[29] <= 32'b011100_00000000000000000000000000; // nop
bios[30] <= 32'b101111_00000_10111_0000000000000000; // rcv $t3
bios[31] <= 32'b010000_11110_10111_1111111111111110; // sw: mem[$sp + (-2)] = mem[$t3]
bios[32] <= 32'b001110_11110_01101_1111111111111110; // lw: $s3 = mem[$sp] + (-2)
bios[33] <= 32'b011011_01101_00110_0000000000000000; // mov: $a0 = $s3
bios[34] <= 32'b111111_00000_00110_0000000000000000; // out $a0
bios[35] <= 32'b001101_11110_11110_0000000000000101; // subi: $sp = $sp - (5)
bios[36] <= 32'b011101_00000000000000000000000000; // hlt*/









		end
	
	always @(posedge clk_auto)
		begin
			biosOut <= bios[address];
		end

	
endmodule

